Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug  9 01:13 2025
                   0fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                   0fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                   2fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                   2fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                   2fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                   2fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                   6fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                   6fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                   6fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                   6fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  10fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  10fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  10fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  10fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  14fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  14fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  14fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  14fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  18fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  18fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  18fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  18fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  22fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  22fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  22fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  22fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  26fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  26fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  26fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  26fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  30fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  30fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  30fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  30fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  34fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  34fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  34fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  34fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  38fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  38fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  38fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  38fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  42fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  42fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  42fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  42fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  46fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  46fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  46fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  46fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  50fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  50fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  50fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  50fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  54fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  54fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  54fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  54fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  58fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  58fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  58fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  58fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  62fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  62fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  62fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  62fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  66fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  66fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  66fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  66fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  70fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  70fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  70fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  70fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  74fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  74fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  74fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                  74fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                  78fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                  78fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                  78fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  78fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                  82fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                  82fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                  82fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  82fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  86fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  86fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  86fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  86fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  90fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                  90fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                  90fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  90fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  94fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  94fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  94fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  94fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                  98fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                  98fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                  98fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                  98fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 102fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 102fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 102fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 102fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 106fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 106fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 106fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 106fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 110fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 110fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 110fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 110fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 114fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 114fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 114fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 114fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 118fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 118fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 118fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 118fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 122fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 122fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 122fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 122fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 126fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 126fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 126fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 126fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 130fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 130fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 130fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 130fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 134fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 134fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 134fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 134fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 138fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 138fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 138fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 138fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 142fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 142fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 142fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 142fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 146fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 146fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 146fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 146fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 150fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 150fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 150fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 150fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 154fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 154fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 154fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 154fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 158fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 158fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 158fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 158fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 162fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 162fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 162fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 162fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 166fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 166fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 166fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 166fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 170fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 170fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 170fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 170fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 174fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 174fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 174fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 174fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 178fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 178fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 178fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 178fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 182fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 182fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 182fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 182fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 186fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 186fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 186fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 186fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 190fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 190fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 190fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 190fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 194fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 194fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 194fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 194fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 198fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 198fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 198fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 198fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 202fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 202fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 202fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 202fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 206fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 206fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 206fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 206fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 210fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 210fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 210fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 210fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 214fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 214fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 214fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 214fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 218fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 218fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 218fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 218fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 222fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 222fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 222fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 222fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 226fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 226fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 226fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 226fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 230fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 230fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 230fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 230fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 234fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 234fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 234fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 234fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 238fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 238fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 238fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 238fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 242fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 242fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 242fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 242fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 246fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 246fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 246fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 246fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 250fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 250fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 250fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 250fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 254fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 254fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 254fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 254fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 258fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 258fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 258fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 258fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 262fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 262fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 262fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 262fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 266fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 266fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 266fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 266fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 270fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 270fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 270fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 270fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 274fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 274fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 274fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 274fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 278fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 278fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 278fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 278fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 282fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 282fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 282fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 282fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 286fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 286fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 286fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 286fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 290fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 290fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 290fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 290fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 294fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 294fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 294fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 294fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 298fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 298fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 298fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 298fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 302fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 302fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 302fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 302fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 306fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 306fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 306fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 306fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 310fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 310fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 310fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 310fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 314fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 314fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 314fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 314fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 318fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 318fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 318fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 318fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 322fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 322fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 322fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 322fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 326fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 326fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 326fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 326fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 330fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 330fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 330fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 330fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 334fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 334fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 334fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 334fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 338fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 338fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 338fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 338fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 342fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 342fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 342fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 342fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 346fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 346fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 346fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 346fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 350fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 350fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 350fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 350fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 354fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 354fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 354fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 354fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 358fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 358fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 358fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 358fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 362fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 362fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 362fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 362fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 366fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 366fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 366fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 366fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 370fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 370fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 370fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 370fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 374fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 374fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 374fr_gen,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 374fr_div,
 rs=1,d_in=0,q_out=0,qb_tog=0
                 378fr_mon,
 rs=1,d_in=0,q_out=0,qb_tog=1
                 378fr_scrb,
 rs=1,d_in=0,q_out=0,qb_tog=1
 done
                 378fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 378fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 382fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 382fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 382fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 382fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 386fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 386fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 386fr_gen,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 386fr_div,
 rs=0,d_in=0,q_out=0,qb_tog=0
                 390fr_mon,
 rs=0,d_in=0,q_out=0,qb_tog=1
                 390fr_scrb,
 rs=0,d_in=0,q_out=0,qb_tog=1
 done
                 390fr_gen,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 390fr_div,
 rs=1,d_in=1,q_out=0,qb_tog=0
                 394fr_mon,
 rs=1,d_in=1,q_out=1,qb_tog=0
                 394fr_scrb,
 rs=1,d_in=1,q_out=1,qb_tog=0
 not_done
                 394fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 394fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 398fr_mon,
 rs=0,d_in=1,q_out=0,qb_tog=1
                 398fr_scrb,
 rs=0,d_in=1,q_out=0,qb_tog=1
 not_done
                 398fr_gen,
 rs=0,d_in=1,q_out=0,qb_tog=0
                 398fr_div,
 rs=0,d_in=1,q_out=0,qb_tog=0
$finish called from file "testbench.sv", line 13.
$finish at simulation time                  400
           V C S   S i m u l a t i o n   R e p o r t 
Time: 400 ns
CPU Time:      0.340 seconds;       Data structure size:   0.0Mb
Sat Aug  9 01:13:20 2025
Done
