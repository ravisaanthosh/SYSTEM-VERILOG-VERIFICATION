interface int_f();
  logic rs,clk;
  logic d_in;
  logic q_out,qb_tog;
endinterface
