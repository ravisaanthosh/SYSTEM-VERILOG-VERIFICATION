interface in_fa;
  logic a;
   logic b;
   logic cin;
   logic sum;
   logic carry;
  endinterface
  
